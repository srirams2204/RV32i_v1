module imm_gen (
    output reg [31:0] imm_out,
    input instr,
    input  [2:0] imm_sel, // 0: I-type, 1: S-type, 2: B-type, 3: U-type, 4: J-type 
);


    
endmodule